--
-- VHDL Architecture fahim_segment_lib.lutled.rtl
--
-- Created:
--          by - user.UNKNOWN (KTP12R7182)
--          at - 13:48:09 01/05/2018
--
-- using Mentor Graphics HDL Designer(TM) 2016.2 (Build 5)
--

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

entity lutled is
  
  port(
    
  d0  : in std_logic_vector(3 downto 0);
  d1  : in std_logic_vector(3 downto 0);
  d2  : in std_logic_vector(3 downto 0);
  d3  : in std_logic_vector(3 downto 0);
 
  spi : out std_logic_vector(31 downto 0)
  
  );
end entity lutled;

--
architecture rtl of lutled is
  signal d0_int           :std_logic_vector(31 downto 0);
  signal d1_int           : std_logic_vector(31 downto 0);
  signal d2_int           : std_logic_vector(31 downto 0);
  signal d3_int           : std_logic_vector(31 downto 0);
 
  
  
begin
  
  with d0 select
  d0_int     <= "00011010111000000000000000000000"   when   "0000",
                "00000010100000000000000000000000"   when   "0001",
                "00011100110000000000000000000000"   when   "0010",
                "00001110110000000000000000000000"   when   "0011",
                "00000110101000000000000000000000"   when   "0100",
                "00001110011000000000000000000000"   when   "0101",
                "00011110011000000000000000000000"   when   "0110",
                "00000010110000000000000000000000"   when   "0111",
                "00011110111000000000000000000000"   when   "1000",
                "00000110111000000000000000000000"   when   "1001",
                "00000000000000000000000000000000"   when   others;

                
  with d1 select              
  d1_int     <= "11000000000110110000000000000000"   when   "0000",
                "01000000000000010000000000000000"   when   "0001",
                "10000000000101110000000000000000"   when   "0010",
                "11000000000001110000000000000000"   when   "0011",
                "01000000000011010000000000000000"   when   "0100",
                "11000000000011100000000000000000"   when   "0101",
                "11000000000111100000000000000000"   when   "0110",
                "01000000000000110000000000000000"   when   "0111",
                "11000000000111110000000000000000"   when   "1000",
                "01000000000011110000000000000000"   when   "1001",
                "00000000000000000000000000000000"   when   others;

                
  with d2 select              
  d2_int     <= "00000000000000000001101011100000"   when   "0000",
                "00000000000000000000001010000000"   when   "0001",
                "00000000000000000001110011000000"   when   "0010",
                "00000000000000000000111011000000"   when   "0011",
                "00000000000000000000011010100000"   when   "0100",
                "00000000000000000000111001100000"   when   "0101",
                "00000000000000000001111001100000"   when   "0110",
                "00000000000000000000001011000000"   when   "0111",
                "00000000000000000001111011100000"   when   "1000",
                "00000000000000000000011011100000"   when   "1001",
                "00000000000000000000000000000000"   when   others;


  with d3 select              
  d3_int     <= "00000000000000001100000000011011"   when   "0000",
                "00000000000000000100000000000001"   when   "0001",
                "00000000000000001000000000010111"   when   "0010",
                "00000000000000001100000000000111"   when   "0011",
                "00000000000000000100000000001101"   when   "0100",
                "00000000000000001100000000001110"   when   "0101",
                "00000000000000001100000000011110"   when   "0110",
                "00000000000000000100000000000011"   when   "0111",
                "00000000000000001100000000011111"   when   "1000",
                "00000000000000000100000000001111"   when   "1001",
                "00000000000000000000000000000000"   when   others;


                
  
  
  spi<= d0_int OR d1_int OR d2_int OR d3_int ;    
        
 
      
end architecture rtl;

